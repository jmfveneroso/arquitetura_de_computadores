library verilog;
use verilog.vl_types.all;
entity Microprocessor is
    port(
        CLK             : in     vl_logic;
        RST             : in     vl_logic
    );
end Microprocessor;
