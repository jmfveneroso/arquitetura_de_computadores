library verilog;
use verilog.vl_types.all;
entity WrapperDE2 is
    port(
        SW15            : in     vl_logic;
        SW14            : in     vl_logic;
        SW13            : in     vl_logic;
        SW12            : in     vl_logic;
        SW11            : in     vl_logic;
        SW10            : in     vl_logic;
        SW9             : in     vl_logic;
        SW8             : in     vl_logic;
        SW7             : in     vl_logic;
        SW6             : in     vl_logic;
        SW5             : in     vl_logic;
        SW4             : in     vl_logic;
        SW3             : in     vl_logic;
        SW2             : in     vl_logic;
        SW1             : in     vl_logic;
        SW0             : in     vl_logic;
        Hex0D0          : out    vl_logic;
        Hex0D1          : out    vl_logic;
        Hex0D2          : out    vl_logic;
        Hex0D3          : out    vl_logic;
        Hex0D4          : out    vl_logic;
        Hex0D5          : out    vl_logic;
        Hex0D6          : out    vl_logic;
        Hex1D0          : out    vl_logic;
        Hex1D1          : out    vl_logic;
        Hex1D2          : out    vl_logic;
        Hex1D3          : out    vl_logic;
        Hex1D4          : out    vl_logic;
        Hex1D5          : out    vl_logic;
        Hex1D6          : out    vl_logic;
        Hex2D0          : out    vl_logic;
        Hex2D1          : out    vl_logic;
        Hex2D2          : out    vl_logic;
        Hex2D3          : out    vl_logic;
        Hex2D4          : out    vl_logic;
        Hex2D5          : out    vl_logic;
        Hex2D6          : out    vl_logic;
        Hex3D0          : out    vl_logic;
        Hex3D1          : out    vl_logic;
        Hex3D2          : out    vl_logic;
        Hex3D3          : out    vl_logic;
        Hex3D4          : out    vl_logic;
        Hex3D5          : out    vl_logic;
        Hex3D6          : out    vl_logic;
        Hex4D0          : out    vl_logic;
        Hex4D1          : out    vl_logic;
        Hex4D2          : out    vl_logic;
        Hex4D3          : out    vl_logic;
        Hex4D4          : out    vl_logic;
        Hex4D5          : out    vl_logic;
        Hex4D6          : out    vl_logic;
        Hex5D0          : out    vl_logic;
        Hex5D1          : out    vl_logic;
        Hex5D2          : out    vl_logic;
        Hex5D3          : out    vl_logic;
        Hex5D4          : out    vl_logic;
        Hex5D5          : out    vl_logic;
        Hex5D6          : out    vl_logic;
        Hex6D0          : out    vl_logic;
        Hex6D1          : out    vl_logic;
        Hex6D2          : out    vl_logic;
        Hex6D3          : out    vl_logic;
        Hex6D4          : out    vl_logic;
        Hex6D5          : out    vl_logic;
        Hex6D6          : out    vl_logic;
        Hex7D0          : out    vl_logic;
        Hex7D1          : out    vl_logic;
        Hex7D2          : out    vl_logic;
        Hex7D3          : out    vl_logic;
        Hex7D4          : out    vl_logic;
        Hex7D5          : out    vl_logic;
        Hex7D6          : out    vl_logic;
        KEY0            : in     vl_logic;
        KEY3            : in     vl_logic;
        CLK             : in     vl_logic;
        RST             : in     vl_logic;
        GO              : in     vl_logic
    );
end WrapperDE2;
