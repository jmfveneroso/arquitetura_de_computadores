library verilog;
use verilog.vl_types.all;
entity Control is
    generic(
        InsADD          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        InsSUB          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        InsSLTI         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        InsAND          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        InsOR           : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        InsXOR          : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        InsANDI         : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi0);
        InsORI          : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        InsXORI         : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        InsADDI         : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi1);
        InsSUBI         : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi0);
        InsJ            : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi1);
        InsBEZ          : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi0);
        InsMUL          : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi0, Hi1);
        InsGHI          : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi0);
        InsGLO          : vl_logic_vector(0 to 3) := (Hi1, Hi1, Hi1, Hi1);
        ULAADD          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        ULASUB          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        ULASLT          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        ULAAND          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        ULAOR           : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        ULAXOR          : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        ULABEZ          : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi0);
        \IF\            : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        ID              : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        RF              : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        EX              : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        WB              : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0)
    );
    port(
        OpCode          : in     vl_logic_vector(3 downto 0);
        ULA_OP          : out    vl_logic_vector(3 downto 0);
        ULA_B           : out    vl_logic;
        EscIR           : out    vl_logic;
        EscCondCP       : out    vl_logic;
        EscCP           : out    vl_logic;
        EscReg          : out    vl_logic;
        WEnPC           : out    vl_logic;
        IsMulWB         : out    vl_logic;
        HILO            : out    vl_logic;
        HILO_WB         : out    vl_logic;
        CLK             : in     vl_logic;
        RST             : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of InsADD : constant is 1;
    attribute mti_svvh_generic_type of InsSUB : constant is 1;
    attribute mti_svvh_generic_type of InsSLTI : constant is 1;
    attribute mti_svvh_generic_type of InsAND : constant is 1;
    attribute mti_svvh_generic_type of InsOR : constant is 1;
    attribute mti_svvh_generic_type of InsXOR : constant is 1;
    attribute mti_svvh_generic_type of InsANDI : constant is 1;
    attribute mti_svvh_generic_type of InsORI : constant is 1;
    attribute mti_svvh_generic_type of InsXORI : constant is 1;
    attribute mti_svvh_generic_type of InsADDI : constant is 1;
    attribute mti_svvh_generic_type of InsSUBI : constant is 1;
    attribute mti_svvh_generic_type of InsJ : constant is 1;
    attribute mti_svvh_generic_type of InsBEZ : constant is 1;
    attribute mti_svvh_generic_type of InsMUL : constant is 1;
    attribute mti_svvh_generic_type of InsGHI : constant is 1;
    attribute mti_svvh_generic_type of InsGLO : constant is 1;
    attribute mti_svvh_generic_type of ULAADD : constant is 1;
    attribute mti_svvh_generic_type of ULASUB : constant is 1;
    attribute mti_svvh_generic_type of ULASLT : constant is 1;
    attribute mti_svvh_generic_type of ULAAND : constant is 1;
    attribute mti_svvh_generic_type of ULAOR : constant is 1;
    attribute mti_svvh_generic_type of ULAXOR : constant is 1;
    attribute mti_svvh_generic_type of ULABEZ : constant is 1;
    attribute mti_svvh_generic_type of \IF\ : constant is 1;
    attribute mti_svvh_generic_type of ID : constant is 1;
    attribute mti_svvh_generic_type of RF : constant is 1;
    attribute mti_svvh_generic_type of EX : constant is 1;
    attribute mti_svvh_generic_type of WB : constant is 1;
end Control;
